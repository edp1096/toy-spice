* BJT Test Circuit
VCC 1 0 DC 10
RB 1 2 100k
Q1 3 2 0 Q2N3904
RC 1 3 1k

.model Q2N3904 NPN(Is=1e-14 Bf=100 Vaf=100)

.tran 1u 1m