* RL Test
.tran 10u 2ms
Vin 1 0 SIN (0 5 1k)
R1 1 2 100
L1 2 0 1m
