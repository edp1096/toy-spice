* Simple BJT AC Test Circuit
VCC 1 0 DC 10
VAC 2 0 AC 0.01
RB 1 2 100k
RC 1 3 10k
Q1 3 2 0 Q2N3904
.model Q2N3904 NPN(Is=1e-14 Bf=100 Vaf=100 Cje=8p Cjc=5p Tf=0.1n Tr=10n)
.ac dec 10 10 1meg