* Simple NMOS Test Circuit

VDD 1 0 DC 5
VG 2 0 PULSE(0 5 1u 100n 100n 5u 10u)

RD 1 3 10k
M1 3 2 0 0 NMOS_Test L=2u W=20u

.model NMOS_Test NMOS(Level=1 VTO=0.7 KP=20u LAMBDA=0.01)

.tran 0.1u 10u
