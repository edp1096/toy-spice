* Transformer Test Circuit with 2:1 ratio
Vin 1 0 sin(0 10 1k)

Rp_leak 1 2 0.1
Lp 2 0 200m

Ls 3 0 50m
Rs_leak 3 4 0.05

Rload 4 0 10k

K1 Lp Ls 0.95

.tran 0.01m 3m