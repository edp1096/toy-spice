* BJT Test Circuit with Base Switching
VCC 1 0 DC 10
VB 4 0 PULSE(0 5 0 1u 1u 100u 200u)
RB 4 2 10
Q1 3 2 0 Q2N3904
RC 1 3 10k

.model Q2N3904 NPN(Is=1e-14 Bf=100 Vaf=100 Cje=10p Cjc=5p Tf=0.3n)
.tran 1u 150u