* RLC Test
.tran 0.1m 3ms
Vin 1 0 SIN(0 5 1k)
R1 1 2 100
L1 2 3 1m
C1 3 0 1u
