* RC Test
.tran 0.01ms 3ms
vin 1 0 sin (0 5 1k)
*.op
*vin 1 0 DC 5
*vin 1 0 ac 1
*.ac dec 10 1 1meg
*.ac lin 100 1 1meg
r1 1 2 100
c1 2 0 1u